`define TEST_MACRO 256
