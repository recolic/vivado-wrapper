`define TEST_MACRO 427