module mod1(
    input i,
    output wire j
);
    assign j = i;
endmodule // mod1